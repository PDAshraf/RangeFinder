-- Range_finder.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity Range_finder is
	port (
		clk_clk            : in  std_logic                    := '0';             --         clk.clk
		distance_in_export : in  std_logic_vector(8 downto 0) := (others => '0'); -- distance_in.export
		ext_irq_export     : in  std_logic_vector(1 downto 0) := (others => '0'); --     ext_irq.export
		key_in_export      : in  std_logic_vector(1 downto 0) := (others => '0'); --      key_in.export
		reset_reset_n      : in  std_logic                    := '0';             --       reset.reset_n
		servo_pos_export   : out std_logic;                                       --   servo_pos.export
		sw_in_export       : in  std_logic_vector(7 downto 0) := (others => '0'); --       sw_in.export
		task_id_export     : out std_logic_vector(2 downto 0);                    --     task_id.export
		vga_b_export       : out std_logic_vector(3 downto 0);                    --       vga_b.export
		vga_g_export       : out std_logic_vector(3 downto 0);                    --       vga_g.export
		vga_hs_export      : out std_logic;                                       --      vga_hs.export
		vga_r_export       : out std_logic_vector(3 downto 0);                    --       vga_r.export
		vga_vs_export      : out std_logic;                                       --      vga_vs.export
		wd_rst_export      : out std_logic                                        --      wd_rst.export
	);
end entity Range_finder;

architecture rtl of Range_finder is
	component SERVO_HW_IP is
		port (
			clk     : in  std_logic                     := 'X';             -- clk
			reset_n : in  std_logic                     := 'X';             -- reset_n
			cs_n    : in  std_logic                     := 'X';             -- chipselect_n
			write_n : in  std_logic                     := 'X';             -- write_n
			din     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			o_pos   : out std_logic                                         -- export
		);
	end component SERVO_HW_IP;

	component TIMER_HW_IP is
		port (
			reset_n : in  std_logic                     := 'X';             -- reset_n
			clk     : in  std_logic                     := 'X';             -- clk
			cs_n    : in  std_logic                     := 'X';             -- chipselect_n
			addr    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n : in  std_logic                     := 'X';             -- write_n
			read_n  : in  std_logic                     := 'X';             -- read_n
			din     : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dout    : out std_logic_vector(31 downto 0)                     -- readdata
		);
	end component TIMER_HW_IP;

	component VGA_IP is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			addr     : in  std_logic_vector(16 downto 0) := (others => 'X'); -- address
			cs_n     : in  std_logic                     := 'X';             -- chipselect_n
			read_n   : in  std_logic                     := 'X';             -- read_n
			write_n  : in  std_logic                     := 'X';             -- write_n
			din      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dout     : out std_logic_vector(31 downto 0);                    -- readdata
			clock_25 : in  std_logic                     := 'X';             -- clk
			vga_r    : out std_logic_vector(3 downto 0);                     -- export
			vga_g    : out std_logic_vector(3 downto 0);                     -- export
			vga_b    : out std_logic_vector(3 downto 0);                     -- export
			vga_hs   : out std_logic;                                        -- export
			vga_vs   : out std_logic                                         -- export
		);
	end component VGA_IP;

	component Range_finder_button_pio is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component Range_finder_button_pio;

	component Range_finder_cpu is
		port (
			clk                                 : in  std_logic                     := 'X';             -- clk
			reset_n                             : in  std_logic                     := 'X';             -- reset_n
			reset_req                           : in  std_logic                     := 'X';             -- reset_req
			d_address                           : out std_logic_vector(19 downto 0);                    -- address
			d_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			d_read                              : out std_logic;                                        -- read
			d_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			d_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			d_write                             : out std_logic;                                        -- write
			d_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			debug_mem_slave_debugaccess_to_roms : out std_logic;                                        -- debugaccess
			i_address                           : out std_logic_vector(19 downto 0);                    -- address
			i_read                              : out std_logic;                                        -- read
			i_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			i_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			irq                                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- irq
			debug_reset_request                 : out std_logic;                                        -- reset
			debug_mem_slave_address             : in  std_logic_vector(8 downto 0)  := (others => 'X'); -- address
			debug_mem_slave_byteenable          : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			debug_mem_slave_debugaccess         : in  std_logic                     := 'X';             -- debugaccess
			debug_mem_slave_read                : in  std_logic                     := 'X';             -- read
			debug_mem_slave_readdata            : out std_logic_vector(31 downto 0);                    -- readdata
			debug_mem_slave_waitrequest         : out std_logic;                                        -- waitrequest
			debug_mem_slave_write               : in  std_logic                     := 'X';             -- write
			debug_mem_slave_writedata           : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			dummy_ci_port                       : out std_logic                                         -- readra
		);
	end component Range_finder_cpu;

	component Range_finder_distance_in is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(8 downto 0)  := (others => 'X')  -- export
		);
	end component Range_finder_distance_in;

	component Range_finder_jtag_uart is
		port (
			clk            : in  std_logic                     := 'X';             -- clk
			rst_n          : in  std_logic                     := 'X';             -- reset_n
			av_chipselect  : in  std_logic                     := 'X';             -- chipselect
			av_address     : in  std_logic                     := 'X';             -- address
			av_read_n      : in  std_logic                     := 'X';             -- read_n
			av_readdata    : out std_logic_vector(31 downto 0);                    -- readdata
			av_write_n     : in  std_logic                     := 'X';             -- write_n
			av_writedata   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			av_waitrequest : out std_logic;                                        -- waitrequest
			av_irq         : out std_logic                                         -- irq
		);
	end component Range_finder_jtag_uart;

	component Range_finder_onchip_ram is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			address    : in  std_logic_vector(14 downto 0) := (others => 'X'); -- address
			clken      : in  std_logic                     := 'X';             -- clken
			chipselect : in  std_logic                     := 'X';             -- chipselect
			write      : in  std_logic                     := 'X';             -- write
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			byteenable : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			reset      : in  std_logic                     := 'X';             -- reset
			reset_req  : in  std_logic                     := 'X';             -- reset_req
			freeze     : in  std_logic                     := 'X'              -- freeze
		);
	end component Range_finder_onchip_ram;

	component Range_finder_pio_out_wd is
		port (
			clk        : in  std_logic                     := 'X';             -- clk
			reset_n    : in  std_logic                     := 'X';             -- reset_n
			address    : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			write_n    : in  std_logic                     := 'X';             -- write_n
			writedata  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			chipselect : in  std_logic                     := 'X';             -- chipselect
			readdata   : out std_logic_vector(31 downto 0);                    -- readdata
			out_port   : out std_logic                                         -- export
		);
	end component Range_finder_pio_out_wd;

	component Range_finder_pll is
		port (
			clk                : in  std_logic                     := 'X';             -- clk
			reset              : in  std_logic                     := 'X';             -- reset
			read               : in  std_logic                     := 'X';             -- read
			write              : in  std_logic                     := 'X';             -- write
			address            : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata           : out std_logic_vector(31 downto 0);                    -- readdata
			writedata          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			c0                 : out std_logic;                                        -- clk
			c1                 : out std_logic;                                        -- clk
			scandone           : out std_logic;                                        -- export
			scandataout        : out std_logic;                                        -- export
			c2                 : out std_logic;                                        -- clk
			c3                 : out std_logic;                                        -- clk
			c4                 : out std_logic;                                        -- clk
			areset             : in  std_logic                     := 'X';             -- export
			locked             : out std_logic;                                        -- export
			phasedone          : out std_logic;                                        -- export
			phasecounterselect : in  std_logic_vector(2 downto 0)  := (others => 'X'); -- export
			phaseupdown        : in  std_logic                     := 'X';             -- export
			phasestep          : in  std_logic                     := 'X';             -- export
			scanclk            : in  std_logic                     := 'X';             -- export
			scanclkena         : in  std_logic                     := 'X';             -- export
			scandata           : in  std_logic                     := 'X';             -- export
			configupdate       : in  std_logic                     := 'X'              -- export
		);
	end component Range_finder_pll;

	component sierra is
		port (
			address                     : in  std_logic_vector(7 downto 0)  := (others => 'X'); -- address
			chipselect_n                : in  std_logic                     := 'X';             -- chipselect_n
			read_n                      : in  std_logic                     := 'X';             -- read_n
			writedata                   : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			write_n                     : in  std_logic                     := 'X';             -- write_n
			readdata                    : out std_logic_vector(31 downto 0);                    -- readdata
			clk                         : in  std_logic                     := 'X';             -- clk
			reset_n                     : in  std_logic                     := 'X';             -- reset_n
			external_runing_taskid_info : out std_logic_vector(2 downto 0);                     -- export
			irq                         : out std_logic;                                        -- irq
			extirq_n                    : in  std_logic_vector(1 downto 0)  := (others => 'X')  -- export
		);
	end component sierra;

	component Range_finder_switch_pio is
		port (
			clk      : in  std_logic                     := 'X';             -- clk
			reset_n  : in  std_logic                     := 'X';             -- reset_n
			address  : in  std_logic_vector(1 downto 0)  := (others => 'X'); -- address
			readdata : out std_logic_vector(31 downto 0);                    -- readdata
			in_port  : in  std_logic_vector(7 downto 0)  := (others => 'X')  -- export
		);
	end component Range_finder_switch_pio;

	component Range_finder_sysid is
		port (
			clock    : in  std_logic                     := 'X'; -- clk
			reset_n  : in  std_logic                     := 'X'; -- reset_n
			readdata : out std_logic_vector(31 downto 0);        -- readdata
			address  : in  std_logic                     := 'X'  -- address
		);
	end component Range_finder_sysid;

	component Range_finder_mm_interconnect_0 is
		port (
			clk_clk_clk                                           : in  std_logic                     := 'X';             -- clk
			pll_c0_clk                                            : in  std_logic                     := 'X';             -- clk
			cpu_reset_reset_bridge_in_reset_reset                 : in  std_logic                     := 'X';             -- reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset : in  std_logic                     := 'X';             -- reset
			cpu_data_master_address                               : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			cpu_data_master_waitrequest                           : out std_logic;                                        -- waitrequest
			cpu_data_master_byteenable                            : in  std_logic_vector(3 downto 0)  := (others => 'X'); -- byteenable
			cpu_data_master_read                                  : in  std_logic                     := 'X';             -- read
			cpu_data_master_readdata                              : out std_logic_vector(31 downto 0);                    -- readdata
			cpu_data_master_write                                 : in  std_logic                     := 'X';             -- write
			cpu_data_master_writedata                             : in  std_logic_vector(31 downto 0) := (others => 'X'); -- writedata
			cpu_data_master_debugaccess                           : in  std_logic                     := 'X';             -- debugaccess
			cpu_instruction_master_address                        : in  std_logic_vector(19 downto 0) := (others => 'X'); -- address
			cpu_instruction_master_waitrequest                    : out std_logic;                                        -- waitrequest
			cpu_instruction_master_read                           : in  std_logic                     := 'X';             -- read
			cpu_instruction_master_readdata                       : out std_logic_vector(31 downto 0);                    -- readdata
			button_pio_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			button_pio_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_address                           : out std_logic_vector(8 downto 0);                     -- address
			cpu_debug_mem_slave_write                             : out std_logic;                                        -- write
			cpu_debug_mem_slave_read                              : out std_logic;                                        -- read
			cpu_debug_mem_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			cpu_debug_mem_slave_writedata                         : out std_logic_vector(31 downto 0);                    -- writedata
			cpu_debug_mem_slave_byteenable                        : out std_logic_vector(3 downto 0);                     -- byteenable
			cpu_debug_mem_slave_waitrequest                       : in  std_logic                     := 'X';             -- waitrequest
			cpu_debug_mem_slave_debugaccess                       : out std_logic;                                        -- debugaccess
			distance_in_s1_address                                : out std_logic_vector(1 downto 0);                     -- address
			distance_in_s1_readdata                               : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_address                   : out std_logic_vector(0 downto 0);                     -- address
			jtag_uart_avalon_jtag_slave_write                     : out std_logic;                                        -- write
			jtag_uart_avalon_jtag_slave_read                      : out std_logic;                                        -- read
			jtag_uart_avalon_jtag_slave_readdata                  : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			jtag_uart_avalon_jtag_slave_writedata                 : out std_logic_vector(31 downto 0);                    -- writedata
			jtag_uart_avalon_jtag_slave_waitrequest               : in  std_logic                     := 'X';             -- waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                : out std_logic;                                        -- chipselect
			onchip_ram_s1_address                                 : out std_logic_vector(14 downto 0);                    -- address
			onchip_ram_s1_write                                   : out std_logic;                                        -- write
			onchip_ram_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			onchip_ram_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			onchip_ram_s1_byteenable                              : out std_logic_vector(3 downto 0);                     -- byteenable
			onchip_ram_s1_chipselect                              : out std_logic;                                        -- chipselect
			onchip_ram_s1_clken                                   : out std_logic;                                        -- clken
			pio_out_wd_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pio_out_wd_s1_write                                   : out std_logic;                                        -- write
			pio_out_wd_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pio_out_wd_s1_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			pio_out_wd_s1_chipselect                              : out std_logic;                                        -- chipselect
			pll_pll_slave_address                                 : out std_logic_vector(1 downto 0);                     -- address
			pll_pll_slave_write                                   : out std_logic;                                        -- write
			pll_pll_slave_read                                    : out std_logic;                                        -- read
			pll_pll_slave_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			pll_pll_slave_writedata                               : out std_logic_vector(31 downto 0);                    -- writedata
			SERVO_HW_IP_0_avalon_slave_0_write                    : out std_logic;                                        -- write
			SERVO_HW_IP_0_avalon_slave_0_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			SERVO_HW_IP_0_avalon_slave_0_chipselect               : out std_logic;                                        -- chipselect
			sierra_0_avalon_slave_0_address                       : out std_logic_vector(7 downto 0);                     -- address
			sierra_0_avalon_slave_0_write                         : out std_logic;                                        -- write
			sierra_0_avalon_slave_0_read                          : out std_logic;                                        -- read
			sierra_0_avalon_slave_0_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sierra_0_avalon_slave_0_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			sierra_0_avalon_slave_0_chipselect                    : out std_logic;                                        -- chipselect
			switch_pio_s1_address                                 : out std_logic_vector(1 downto 0);                     -- address
			switch_pio_s1_readdata                                : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			sysid_control_slave_address                           : out std_logic_vector(0 downto 0);                     -- address
			sysid_control_slave_readdata                          : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TIMER_HW_IP_0_avalon_slave_0_address                  : out std_logic_vector(1 downto 0);                     -- address
			TIMER_HW_IP_0_avalon_slave_0_write                    : out std_logic;                                        -- write
			TIMER_HW_IP_0_avalon_slave_0_read                     : out std_logic;                                        -- read
			TIMER_HW_IP_0_avalon_slave_0_readdata                 : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			TIMER_HW_IP_0_avalon_slave_0_writedata                : out std_logic_vector(31 downto 0);                    -- writedata
			TIMER_HW_IP_0_avalon_slave_0_chipselect               : out std_logic;                                        -- chipselect
			VGA_IP_0_avalon_slave_0_address                       : out std_logic_vector(16 downto 0);                    -- address
			VGA_IP_0_avalon_slave_0_write                         : out std_logic;                                        -- write
			VGA_IP_0_avalon_slave_0_read                          : out std_logic;                                        -- read
			VGA_IP_0_avalon_slave_0_readdata                      : in  std_logic_vector(31 downto 0) := (others => 'X'); -- readdata
			VGA_IP_0_avalon_slave_0_writedata                     : out std_logic_vector(31 downto 0);                    -- writedata
			VGA_IP_0_avalon_slave_0_chipselect                    : out std_logic                                         -- chipselect
		);
	end component Range_finder_mm_interconnect_0;

	component Range_finder_irq_mapper is
		port (
			clk           : in  std_logic                     := 'X'; -- clk
			reset         : in  std_logic                     := 'X'; -- reset
			receiver0_irq : in  std_logic                     := 'X'; -- irq
			receiver1_irq : in  std_logic                     := 'X'; -- irq
			sender_irq    : out std_logic_vector(31 downto 0)         -- irq
		);
	end component Range_finder_irq_mapper;

	component range_finder_rst_controller is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_req      : out std_logic;        --          .reset_req
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component range_finder_rst_controller;

	component range_finder_rst_controller_001 is
		generic (
			NUM_RESET_INPUTS          : integer := 6;
			OUTPUT_RESET_SYNC_EDGES   : string  := "deassert";
			SYNC_DEPTH                : integer := 2;
			RESET_REQUEST_PRESENT     : integer := 0;
			RESET_REQ_WAIT_TIME       : integer := 1;
			MIN_RST_ASSERTION_TIME    : integer := 3;
			RESET_REQ_EARLY_DSRT_TIME : integer := 1;
			USE_RESET_REQUEST_IN0     : integer := 0;
			USE_RESET_REQUEST_IN1     : integer := 0;
			USE_RESET_REQUEST_IN2     : integer := 0;
			USE_RESET_REQUEST_IN3     : integer := 0;
			USE_RESET_REQUEST_IN4     : integer := 0;
			USE_RESET_REQUEST_IN5     : integer := 0;
			USE_RESET_REQUEST_IN6     : integer := 0;
			USE_RESET_REQUEST_IN7     : integer := 0;
			USE_RESET_REQUEST_IN8     : integer := 0;
			USE_RESET_REQUEST_IN9     : integer := 0;
			USE_RESET_REQUEST_IN10    : integer := 0;
			USE_RESET_REQUEST_IN11    : integer := 0;
			USE_RESET_REQUEST_IN12    : integer := 0;
			USE_RESET_REQUEST_IN13    : integer := 0;
			USE_RESET_REQUEST_IN14    : integer := 0;
			USE_RESET_REQUEST_IN15    : integer := 0;
			ADAPT_RESET_REQUEST       : integer := 0
		);
		port (
			reset_in0      : in  std_logic := 'X'; -- reset_in0.reset
			reset_in1      : in  std_logic := 'X'; -- reset_in1.reset
			clk            : in  std_logic := 'X'; --       clk.clk
			reset_out      : out std_logic;        -- reset_out.reset
			reset_in10     : in  std_logic := 'X';
			reset_in11     : in  std_logic := 'X';
			reset_in12     : in  std_logic := 'X';
			reset_in13     : in  std_logic := 'X';
			reset_in14     : in  std_logic := 'X';
			reset_in15     : in  std_logic := 'X';
			reset_in2      : in  std_logic := 'X';
			reset_in3      : in  std_logic := 'X';
			reset_in4      : in  std_logic := 'X';
			reset_in5      : in  std_logic := 'X';
			reset_in6      : in  std_logic := 'X';
			reset_in7      : in  std_logic := 'X';
			reset_in8      : in  std_logic := 'X';
			reset_in9      : in  std_logic := 'X';
			reset_req      : out std_logic;
			reset_req_in0  : in  std_logic := 'X';
			reset_req_in1  : in  std_logic := 'X';
			reset_req_in10 : in  std_logic := 'X';
			reset_req_in11 : in  std_logic := 'X';
			reset_req_in12 : in  std_logic := 'X';
			reset_req_in13 : in  std_logic := 'X';
			reset_req_in14 : in  std_logic := 'X';
			reset_req_in15 : in  std_logic := 'X';
			reset_req_in2  : in  std_logic := 'X';
			reset_req_in3  : in  std_logic := 'X';
			reset_req_in4  : in  std_logic := 'X';
			reset_req_in5  : in  std_logic := 'X';
			reset_req_in6  : in  std_logic := 'X';
			reset_req_in7  : in  std_logic := 'X';
			reset_req_in8  : in  std_logic := 'X';
			reset_req_in9  : in  std_logic := 'X'
		);
	end component range_finder_rst_controller_001;

	signal pll_c0_clk                                                          : std_logic;                     -- pll:c0 -> [SERVO_HW_IP_0:clk, TIMER_HW_IP_0:clk, VGA_IP_0:clk, button_pio:clk, cpu:clk, distance_in:clk, irq_mapper:clk, jtag_uart:clk, mm_interconnect_0:pll_c0_clk, onchip_ram:clk, pio_out_wd:clk, rst_controller:clk, sierra_0:clk, switch_pio:clk, sysid:clock]
	signal pll_c1_clk                                                          : std_logic;                     -- pll:c1 -> VGA_IP_0:clock_25
	signal cpu_data_master_readdata                                            : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_data_master_readdata -> cpu:d_readdata
	signal cpu_data_master_waitrequest                                         : std_logic;                     -- mm_interconnect_0:cpu_data_master_waitrequest -> cpu:d_waitrequest
	signal cpu_data_master_debugaccess                                         : std_logic;                     -- cpu:debug_mem_slave_debugaccess_to_roms -> mm_interconnect_0:cpu_data_master_debugaccess
	signal cpu_data_master_address                                             : std_logic_vector(19 downto 0); -- cpu:d_address -> mm_interconnect_0:cpu_data_master_address
	signal cpu_data_master_byteenable                                          : std_logic_vector(3 downto 0);  -- cpu:d_byteenable -> mm_interconnect_0:cpu_data_master_byteenable
	signal cpu_data_master_read                                                : std_logic;                     -- cpu:d_read -> mm_interconnect_0:cpu_data_master_read
	signal cpu_data_master_write                                               : std_logic;                     -- cpu:d_write -> mm_interconnect_0:cpu_data_master_write
	signal cpu_data_master_writedata                                           : std_logic_vector(31 downto 0); -- cpu:d_writedata -> mm_interconnect_0:cpu_data_master_writedata
	signal cpu_instruction_master_readdata                                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_instruction_master_readdata -> cpu:i_readdata
	signal cpu_instruction_master_waitrequest                                  : std_logic;                     -- mm_interconnect_0:cpu_instruction_master_waitrequest -> cpu:i_waitrequest
	signal cpu_instruction_master_address                                      : std_logic_vector(19 downto 0); -- cpu:i_address -> mm_interconnect_0:cpu_instruction_master_address
	signal cpu_instruction_master_read                                         : std_logic;                     -- cpu:i_read -> mm_interconnect_0:cpu_instruction_master_read
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect            : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_chipselect -> jtag_uart:av_chipselect
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata              : std_logic_vector(31 downto 0); -- jtag_uart:av_readdata -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_readdata
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest           : std_logic;                     -- jtag_uart:av_waitrequest -> mm_interconnect_0:jtag_uart_avalon_jtag_slave_waitrequest
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_address               : std_logic_vector(0 downto 0);  -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_address -> jtag_uart:av_address
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read                  : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_read -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write                 : std_logic;                     -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_write -> mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:in
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata             : std_logic_vector(31 downto 0); -- mm_interconnect_0:jtag_uart_avalon_jtag_slave_writedata -> jtag_uart:av_writedata
	signal mm_interconnect_0_sierra_0_avalon_slave_0_chipselect                : std_logic;                     -- mm_interconnect_0:sierra_0_avalon_slave_0_chipselect -> mm_interconnect_0_sierra_0_avalon_slave_0_chipselect:in
	signal mm_interconnect_0_sierra_0_avalon_slave_0_readdata                  : std_logic_vector(31 downto 0); -- sierra_0:readdata -> mm_interconnect_0:sierra_0_avalon_slave_0_readdata
	signal mm_interconnect_0_sierra_0_avalon_slave_0_address                   : std_logic_vector(7 downto 0);  -- mm_interconnect_0:sierra_0_avalon_slave_0_address -> sierra_0:address
	signal mm_interconnect_0_sierra_0_avalon_slave_0_read                      : std_logic;                     -- mm_interconnect_0:sierra_0_avalon_slave_0_read -> mm_interconnect_0_sierra_0_avalon_slave_0_read:in
	signal mm_interconnect_0_sierra_0_avalon_slave_0_write                     : std_logic;                     -- mm_interconnect_0:sierra_0_avalon_slave_0_write -> mm_interconnect_0_sierra_0_avalon_slave_0_write:in
	signal mm_interconnect_0_sierra_0_avalon_slave_0_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:sierra_0_avalon_slave_0_writedata -> sierra_0:writedata
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect                : std_logic;                     -- mm_interconnect_0:VGA_IP_0_avalon_slave_0_chipselect -> mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect:in
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_readdata                  : std_logic_vector(31 downto 0); -- VGA_IP_0:dout -> mm_interconnect_0:VGA_IP_0_avalon_slave_0_readdata
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_address                   : std_logic_vector(16 downto 0); -- mm_interconnect_0:VGA_IP_0_avalon_slave_0_address -> VGA_IP_0:addr
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_read                      : std_logic;                     -- mm_interconnect_0:VGA_IP_0_avalon_slave_0_read -> mm_interconnect_0_vga_ip_0_avalon_slave_0_read:in
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_write                     : std_logic;                     -- mm_interconnect_0:VGA_IP_0_avalon_slave_0_write -> mm_interconnect_0_vga_ip_0_avalon_slave_0_write:in
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_writedata                 : std_logic_vector(31 downto 0); -- mm_interconnect_0:VGA_IP_0_avalon_slave_0_writedata -> VGA_IP_0:din
	signal mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_chipselect           : std_logic;                     -- mm_interconnect_0:SERVO_HW_IP_0_avalon_slave_0_chipselect -> mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_chipselect:in
	signal mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_write                : std_logic;                     -- mm_interconnect_0:SERVO_HW_IP_0_avalon_slave_0_write -> mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_write:in
	signal mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:SERVO_HW_IP_0_avalon_slave_0_writedata -> SERVO_HW_IP_0:din
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect           : std_logic;                     -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_chipselect -> mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect:in
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_readdata             : std_logic_vector(31 downto 0); -- TIMER_HW_IP_0:dout -> mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_readdata
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_address              : std_logic_vector(1 downto 0);  -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_address -> TIMER_HW_IP_0:addr
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read                 : std_logic;                     -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_read -> mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read:in
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write                : std_logic;                     -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_write -> mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write:in
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_writedata            : std_logic_vector(31 downto 0); -- mm_interconnect_0:TIMER_HW_IP_0_avalon_slave_0_writedata -> TIMER_HW_IP_0:din
	signal mm_interconnect_0_sysid_control_slave_readdata                      : std_logic_vector(31 downto 0); -- sysid:readdata -> mm_interconnect_0:sysid_control_slave_readdata
	signal mm_interconnect_0_sysid_control_slave_address                       : std_logic_vector(0 downto 0);  -- mm_interconnect_0:sysid_control_slave_address -> sysid:address
	signal mm_interconnect_0_cpu_debug_mem_slave_readdata                      : std_logic_vector(31 downto 0); -- cpu:debug_mem_slave_readdata -> mm_interconnect_0:cpu_debug_mem_slave_readdata
	signal mm_interconnect_0_cpu_debug_mem_slave_waitrequest                   : std_logic;                     -- cpu:debug_mem_slave_waitrequest -> mm_interconnect_0:cpu_debug_mem_slave_waitrequest
	signal mm_interconnect_0_cpu_debug_mem_slave_debugaccess                   : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_debugaccess -> cpu:debug_mem_slave_debugaccess
	signal mm_interconnect_0_cpu_debug_mem_slave_address                       : std_logic_vector(8 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_address -> cpu:debug_mem_slave_address
	signal mm_interconnect_0_cpu_debug_mem_slave_read                          : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_read -> cpu:debug_mem_slave_read
	signal mm_interconnect_0_cpu_debug_mem_slave_byteenable                    : std_logic_vector(3 downto 0);  -- mm_interconnect_0:cpu_debug_mem_slave_byteenable -> cpu:debug_mem_slave_byteenable
	signal mm_interconnect_0_cpu_debug_mem_slave_write                         : std_logic;                     -- mm_interconnect_0:cpu_debug_mem_slave_write -> cpu:debug_mem_slave_write
	signal mm_interconnect_0_cpu_debug_mem_slave_writedata                     : std_logic_vector(31 downto 0); -- mm_interconnect_0:cpu_debug_mem_slave_writedata -> cpu:debug_mem_slave_writedata
	signal mm_interconnect_0_pll_pll_slave_readdata                            : std_logic_vector(31 downto 0); -- pll:readdata -> mm_interconnect_0:pll_pll_slave_readdata
	signal mm_interconnect_0_pll_pll_slave_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pll_pll_slave_address -> pll:address
	signal mm_interconnect_0_pll_pll_slave_read                                : std_logic;                     -- mm_interconnect_0:pll_pll_slave_read -> pll:read
	signal mm_interconnect_0_pll_pll_slave_write                               : std_logic;                     -- mm_interconnect_0:pll_pll_slave_write -> pll:write
	signal mm_interconnect_0_pll_pll_slave_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:pll_pll_slave_writedata -> pll:writedata
	signal mm_interconnect_0_onchip_ram_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_chipselect -> onchip_ram:chipselect
	signal mm_interconnect_0_onchip_ram_s1_readdata                            : std_logic_vector(31 downto 0); -- onchip_ram:readdata -> mm_interconnect_0:onchip_ram_s1_readdata
	signal mm_interconnect_0_onchip_ram_s1_address                             : std_logic_vector(14 downto 0); -- mm_interconnect_0:onchip_ram_s1_address -> onchip_ram:address
	signal mm_interconnect_0_onchip_ram_s1_byteenable                          : std_logic_vector(3 downto 0);  -- mm_interconnect_0:onchip_ram_s1_byteenable -> onchip_ram:byteenable
	signal mm_interconnect_0_onchip_ram_s1_write                               : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_write -> onchip_ram:write
	signal mm_interconnect_0_onchip_ram_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:onchip_ram_s1_writedata -> onchip_ram:writedata
	signal mm_interconnect_0_onchip_ram_s1_clken                               : std_logic;                     -- mm_interconnect_0:onchip_ram_s1_clken -> onchip_ram:clken
	signal mm_interconnect_0_distance_in_s1_readdata                           : std_logic_vector(31 downto 0); -- distance_in:readdata -> mm_interconnect_0:distance_in_s1_readdata
	signal mm_interconnect_0_distance_in_s1_address                            : std_logic_vector(1 downto 0);  -- mm_interconnect_0:distance_in_s1_address -> distance_in:address
	signal mm_interconnect_0_pio_out_wd_s1_chipselect                          : std_logic;                     -- mm_interconnect_0:pio_out_wd_s1_chipselect -> pio_out_wd:chipselect
	signal mm_interconnect_0_pio_out_wd_s1_readdata                            : std_logic_vector(31 downto 0); -- pio_out_wd:readdata -> mm_interconnect_0:pio_out_wd_s1_readdata
	signal mm_interconnect_0_pio_out_wd_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:pio_out_wd_s1_address -> pio_out_wd:address
	signal mm_interconnect_0_pio_out_wd_s1_write                               : std_logic;                     -- mm_interconnect_0:pio_out_wd_s1_write -> mm_interconnect_0_pio_out_wd_s1_write:in
	signal mm_interconnect_0_pio_out_wd_s1_writedata                           : std_logic_vector(31 downto 0); -- mm_interconnect_0:pio_out_wd_s1_writedata -> pio_out_wd:writedata
	signal mm_interconnect_0_button_pio_s1_readdata                            : std_logic_vector(31 downto 0); -- button_pio:readdata -> mm_interconnect_0:button_pio_s1_readdata
	signal mm_interconnect_0_button_pio_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:button_pio_s1_address -> button_pio:address
	signal mm_interconnect_0_switch_pio_s1_readdata                            : std_logic_vector(31 downto 0); -- switch_pio:readdata -> mm_interconnect_0:switch_pio_s1_readdata
	signal mm_interconnect_0_switch_pio_s1_address                             : std_logic_vector(1 downto 0);  -- mm_interconnect_0:switch_pio_s1_address -> switch_pio:address
	signal irq_mapper_receiver0_irq                                            : std_logic;                     -- sierra_0:irq -> irq_mapper:receiver0_irq
	signal irq_mapper_receiver1_irq                                            : std_logic;                     -- jtag_uart:av_irq -> irq_mapper:receiver1_irq
	signal cpu_irq_irq                                                         : std_logic_vector(31 downto 0); -- irq_mapper:sender_irq -> cpu:irq
	signal rst_controller_reset_out_reset                                      : std_logic;                     -- rst_controller:reset_out -> [irq_mapper:reset, mm_interconnect_0:cpu_reset_reset_bridge_in_reset_reset, onchip_ram:reset, rst_controller_reset_out_reset:in, rst_translator:in_reset]
	signal rst_controller_reset_out_reset_req                                  : std_logic;                     -- rst_controller:reset_req -> [cpu:reset_req, onchip_ram:reset_req, rst_translator:reset_req_in]
	signal cpu_debug_reset_request_reset                                       : std_logic;                     -- cpu:debug_reset_request -> [rst_controller:reset_in1, rst_controller_001:reset_in1]
	signal rst_controller_001_reset_out_reset                                  : std_logic;                     -- rst_controller_001:reset_out -> [mm_interconnect_0:pll_inclk_interface_reset_reset_bridge_in_reset_reset, pll:reset]
	signal reset_reset_n_ports_inv                                             : std_logic;                     -- reset_reset_n:inv -> [rst_controller:reset_in0, rst_controller_001:reset_in0]
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv        : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_read:inv -> jtag_uart:av_read_n
	signal mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv       : std_logic;                     -- mm_interconnect_0_jtag_uart_avalon_jtag_slave_write:inv -> jtag_uart:av_write_n
	signal mm_interconnect_0_sierra_0_avalon_slave_0_chipselect_ports_inv      : std_logic;                     -- mm_interconnect_0_sierra_0_avalon_slave_0_chipselect:inv -> sierra_0:chipselect_n
	signal mm_interconnect_0_sierra_0_avalon_slave_0_read_ports_inv            : std_logic;                     -- mm_interconnect_0_sierra_0_avalon_slave_0_read:inv -> sierra_0:read_n
	signal mm_interconnect_0_sierra_0_avalon_slave_0_write_ports_inv           : std_logic;                     -- mm_interconnect_0_sierra_0_avalon_slave_0_write:inv -> sierra_0:write_n
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect_ports_inv      : std_logic;                     -- mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect:inv -> VGA_IP_0:cs_n
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_read_ports_inv            : std_logic;                     -- mm_interconnect_0_vga_ip_0_avalon_slave_0_read:inv -> VGA_IP_0:read_n
	signal mm_interconnect_0_vga_ip_0_avalon_slave_0_write_ports_inv           : std_logic;                     -- mm_interconnect_0_vga_ip_0_avalon_slave_0_write:inv -> VGA_IP_0:write_n
	signal mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_chipselect_ports_inv : std_logic;                     -- mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_chipselect:inv -> SERVO_HW_IP_0:cs_n
	signal mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_write_ports_inv      : std_logic;                     -- mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_write:inv -> SERVO_HW_IP_0:write_n
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect_ports_inv : std_logic;                     -- mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect:inv -> TIMER_HW_IP_0:cs_n
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read_ports_inv       : std_logic;                     -- mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read:inv -> TIMER_HW_IP_0:read_n
	signal mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write_ports_inv      : std_logic;                     -- mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write:inv -> TIMER_HW_IP_0:write_n
	signal mm_interconnect_0_pio_out_wd_s1_write_ports_inv                     : std_logic;                     -- mm_interconnect_0_pio_out_wd_s1_write:inv -> pio_out_wd:write_n
	signal rst_controller_reset_out_reset_ports_inv                            : std_logic;                     -- rst_controller_reset_out_reset:inv -> [SERVO_HW_IP_0:reset_n, TIMER_HW_IP_0:reset_n, VGA_IP_0:reset_n, button_pio:reset_n, cpu:reset_n, distance_in:reset_n, jtag_uart:rst_n, pio_out_wd:reset_n, sierra_0:reset_n, switch_pio:reset_n, sysid:reset_n]

begin

	servo_hw_ip_0 : component SERVO_HW_IP
		port map (
			clk     => pll_c0_clk,                                                          --          clock.clk
			reset_n => rst_controller_reset_out_reset_ports_inv,                            --          reset.reset_n
			cs_n    => mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_chipselect_ports_inv, -- avalon_slave_0.chipselect_n
			write_n => mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_write_ports_inv,      --               .write_n
			din     => mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_writedata,            --               .writedata
			o_pos   => servo_pos_export                                                     --    conduit_end.export
		);

	timer_hw_ip_0 : component TIMER_HW_IP
		port map (
			reset_n => rst_controller_reset_out_reset_ports_inv,                            --          reset.reset_n
			clk     => pll_c0_clk,                                                          --          clock.clk
			cs_n    => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect_ports_inv, -- avalon_slave_0.chipselect_n
			addr    => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_address,              --               .address
			write_n => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write_ports_inv,      --               .write_n
			read_n  => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read_ports_inv,       --               .read_n
			din     => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_writedata,            --               .writedata
			dout    => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_readdata              --               .readdata
		);

	vga_ip_0 : component VGA_IP
		port map (
			clk      => pll_c0_clk,                                                     --          clock.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,                       --          reset.reset_n
			addr     => mm_interconnect_0_vga_ip_0_avalon_slave_0_address,              -- avalon_slave_0.address
			cs_n     => mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect_ports_inv, --               .chipselect_n
			read_n   => mm_interconnect_0_vga_ip_0_avalon_slave_0_read_ports_inv,       --               .read_n
			write_n  => mm_interconnect_0_vga_ip_0_avalon_slave_0_write_ports_inv,      --               .write_n
			din      => mm_interconnect_0_vga_ip_0_avalon_slave_0_writedata,            --               .writedata
			dout     => mm_interconnect_0_vga_ip_0_avalon_slave_0_readdata,             --               .readdata
			clock_25 => pll_c1_clk,                                                     --     clock_sink.clk
			vga_r    => vga_r_export,                                                   --  conduit_end_1.export
			vga_g    => vga_g_export,                                                   --  conduit_end_2.export
			vga_b    => vga_b_export,                                                   --  conduit_end_3.export
			vga_hs   => vga_hs_export,                                                  --  conduit_end_4.export
			vga_vs   => vga_vs_export                                                   --  conduit_end_5.export
		);

	button_pio : component Range_finder_button_pio
		port map (
			clk      => pll_c0_clk,                               --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_button_pio_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_button_pio_s1_readdata, --                    .readdata
			in_port  => key_in_export                             -- external_connection.export
		);

	cpu : component Range_finder_cpu
		port map (
			clk                                 => pll_c0_clk,                                        --                       clk.clk
			reset_n                             => rst_controller_reset_out_reset_ports_inv,          --                     reset.reset_n
			reset_req                           => rst_controller_reset_out_reset_req,                --                          .reset_req
			d_address                           => cpu_data_master_address,                           --               data_master.address
			d_byteenable                        => cpu_data_master_byteenable,                        --                          .byteenable
			d_read                              => cpu_data_master_read,                              --                          .read
			d_readdata                          => cpu_data_master_readdata,                          --                          .readdata
			d_waitrequest                       => cpu_data_master_waitrequest,                       --                          .waitrequest
			d_write                             => cpu_data_master_write,                             --                          .write
			d_writedata                         => cpu_data_master_writedata,                         --                          .writedata
			debug_mem_slave_debugaccess_to_roms => cpu_data_master_debugaccess,                       --                          .debugaccess
			i_address                           => cpu_instruction_master_address,                    --        instruction_master.address
			i_read                              => cpu_instruction_master_read,                       --                          .read
			i_readdata                          => cpu_instruction_master_readdata,                   --                          .readdata
			i_waitrequest                       => cpu_instruction_master_waitrequest,                --                          .waitrequest
			irq                                 => cpu_irq_irq,                                       --                       irq.irq
			debug_reset_request                 => cpu_debug_reset_request_reset,                     --       debug_reset_request.reset
			debug_mem_slave_address             => mm_interconnect_0_cpu_debug_mem_slave_address,     --           debug_mem_slave.address
			debug_mem_slave_byteenable          => mm_interconnect_0_cpu_debug_mem_slave_byteenable,  --                          .byteenable
			debug_mem_slave_debugaccess         => mm_interconnect_0_cpu_debug_mem_slave_debugaccess, --                          .debugaccess
			debug_mem_slave_read                => mm_interconnect_0_cpu_debug_mem_slave_read,        --                          .read
			debug_mem_slave_readdata            => mm_interconnect_0_cpu_debug_mem_slave_readdata,    --                          .readdata
			debug_mem_slave_waitrequest         => mm_interconnect_0_cpu_debug_mem_slave_waitrequest, --                          .waitrequest
			debug_mem_slave_write               => mm_interconnect_0_cpu_debug_mem_slave_write,       --                          .write
			debug_mem_slave_writedata           => mm_interconnect_0_cpu_debug_mem_slave_writedata,   --                          .writedata
			dummy_ci_port                       => open                                               -- custom_instruction_master.readra
		);

	distance_in : component Range_finder_distance_in
		port map (
			clk      => pll_c0_clk,                                --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,  --               reset.reset_n
			address  => mm_interconnect_0_distance_in_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_distance_in_s1_readdata, --                    .readdata
			in_port  => distance_in_export                         -- external_connection.export
		);

	jtag_uart : component Range_finder_jtag_uart
		port map (
			clk            => pll_c0_clk,                                                    --               clk.clk
			rst_n          => rst_controller_reset_out_reset_ports_inv,                      --             reset.reset_n
			av_chipselect  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,      -- avalon_jtag_slave.chipselect
			av_address     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address(0),      --                  .address
			av_read_n      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv,  --                  .read_n
			av_readdata    => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,        --                  .readdata
			av_write_n     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv, --                  .write_n
			av_writedata   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,       --                  .writedata
			av_waitrequest => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest,     --                  .waitrequest
			av_irq         => irq_mapper_receiver1_irq                                       --               irq.irq
		);

	onchip_ram : component Range_finder_onchip_ram
		port map (
			clk        => pll_c0_clk,                                 --   clk1.clk
			address    => mm_interconnect_0_onchip_ram_s1_address,    --     s1.address
			clken      => mm_interconnect_0_onchip_ram_s1_clken,      --       .clken
			chipselect => mm_interconnect_0_onchip_ram_s1_chipselect, --       .chipselect
			write      => mm_interconnect_0_onchip_ram_s1_write,      --       .write
			readdata   => mm_interconnect_0_onchip_ram_s1_readdata,   --       .readdata
			writedata  => mm_interconnect_0_onchip_ram_s1_writedata,  --       .writedata
			byteenable => mm_interconnect_0_onchip_ram_s1_byteenable, --       .byteenable
			reset      => rst_controller_reset_out_reset,             -- reset1.reset
			reset_req  => rst_controller_reset_out_reset_req,         --       .reset_req
			freeze     => '0'                                         -- (terminated)
		);

	pio_out_wd : component Range_finder_pio_out_wd
		port map (
			clk        => pll_c0_clk,                                      --                 clk.clk
			reset_n    => rst_controller_reset_out_reset_ports_inv,        --               reset.reset_n
			address    => mm_interconnect_0_pio_out_wd_s1_address,         --                  s1.address
			write_n    => mm_interconnect_0_pio_out_wd_s1_write_ports_inv, --                    .write_n
			writedata  => mm_interconnect_0_pio_out_wd_s1_writedata,       --                    .writedata
			chipselect => mm_interconnect_0_pio_out_wd_s1_chipselect,      --                    .chipselect
			readdata   => mm_interconnect_0_pio_out_wd_s1_readdata,        --                    .readdata
			out_port   => wd_rst_export                                    -- external_connection.export
		);

	pll : component Range_finder_pll
		port map (
			clk                => clk_clk,                                   --       inclk_interface.clk
			reset              => rst_controller_001_reset_out_reset,        -- inclk_interface_reset.reset
			read               => mm_interconnect_0_pll_pll_slave_read,      --             pll_slave.read
			write              => mm_interconnect_0_pll_pll_slave_write,     --                      .write
			address            => mm_interconnect_0_pll_pll_slave_address,   --                      .address
			readdata           => mm_interconnect_0_pll_pll_slave_readdata,  --                      .readdata
			writedata          => mm_interconnect_0_pll_pll_slave_writedata, --                      .writedata
			c0                 => pll_c0_clk,                                --                    c0.clk
			c1                 => pll_c1_clk,                                --                    c1.clk
			scandone           => open,                                      --           (terminated)
			scandataout        => open,                                      --           (terminated)
			c2                 => open,                                      --           (terminated)
			c3                 => open,                                      --           (terminated)
			c4                 => open,                                      --           (terminated)
			areset             => '0',                                       --           (terminated)
			locked             => open,                                      --           (terminated)
			phasedone          => open,                                      --           (terminated)
			phasecounterselect => "000",                                     --           (terminated)
			phaseupdown        => '0',                                       --           (terminated)
			phasestep          => '0',                                       --           (terminated)
			scanclk            => '0',                                       --           (terminated)
			scanclkena         => '0',                                       --           (terminated)
			scandata           => '0',                                       --           (terminated)
			configupdate       => '0'                                        --           (terminated)
		);

	sierra_0 : component sierra
		port map (
			address                     => mm_interconnect_0_sierra_0_avalon_slave_0_address,              --    avalon_slave_0.address
			chipselect_n                => mm_interconnect_0_sierra_0_avalon_slave_0_chipselect_ports_inv, --                  .chipselect_n
			read_n                      => mm_interconnect_0_sierra_0_avalon_slave_0_read_ports_inv,       --                  .read_n
			writedata                   => mm_interconnect_0_sierra_0_avalon_slave_0_writedata,            --                  .writedata
			write_n                     => mm_interconnect_0_sierra_0_avalon_slave_0_write_ports_inv,      --                  .write_n
			readdata                    => mm_interconnect_0_sierra_0_avalon_slave_0_readdata,             --                  .readdata
			clk                         => pll_c0_clk,                                                     --       clock_reset.clk
			reset_n                     => rst_controller_reset_out_reset_ports_inv,                       -- clock_reset_reset.reset_n
			external_runing_taskid_info => task_id_export,                                                 --       conduit_end.export
			irq                         => irq_mapper_receiver0_irq,                                       --  interrupt_sender.irq
			extirq_n                    => ext_irq_export                                                  --     conduit_end_1.export
		);

	switch_pio : component Range_finder_switch_pio
		port map (
			clk      => pll_c0_clk,                               --                 clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv, --               reset.reset_n
			address  => mm_interconnect_0_switch_pio_s1_address,  --                  s1.address
			readdata => mm_interconnect_0_switch_pio_s1_readdata, --                    .readdata
			in_port  => sw_in_export                              -- external_connection.export
		);

	sysid : component Range_finder_sysid
		port map (
			clock    => pll_c0_clk,                                       --           clk.clk
			reset_n  => rst_controller_reset_out_reset_ports_inv,         --         reset.reset_n
			readdata => mm_interconnect_0_sysid_control_slave_readdata,   -- control_slave.readdata
			address  => mm_interconnect_0_sysid_control_slave_address(0)  --              .address
		);

	mm_interconnect_0 : component Range_finder_mm_interconnect_0
		port map (
			clk_clk_clk                                           => clk_clk,                                                   --                                         clk_clk.clk
			pll_c0_clk                                            => pll_c0_clk,                                                --                                          pll_c0.clk
			cpu_reset_reset_bridge_in_reset_reset                 => rst_controller_reset_out_reset,                            --                 cpu_reset_reset_bridge_in_reset.reset
			pll_inclk_interface_reset_reset_bridge_in_reset_reset => rst_controller_001_reset_out_reset,                        -- pll_inclk_interface_reset_reset_bridge_in_reset.reset
			cpu_data_master_address                               => cpu_data_master_address,                                   --                                 cpu_data_master.address
			cpu_data_master_waitrequest                           => cpu_data_master_waitrequest,                               --                                                .waitrequest
			cpu_data_master_byteenable                            => cpu_data_master_byteenable,                                --                                                .byteenable
			cpu_data_master_read                                  => cpu_data_master_read,                                      --                                                .read
			cpu_data_master_readdata                              => cpu_data_master_readdata,                                  --                                                .readdata
			cpu_data_master_write                                 => cpu_data_master_write,                                     --                                                .write
			cpu_data_master_writedata                             => cpu_data_master_writedata,                                 --                                                .writedata
			cpu_data_master_debugaccess                           => cpu_data_master_debugaccess,                               --                                                .debugaccess
			cpu_instruction_master_address                        => cpu_instruction_master_address,                            --                          cpu_instruction_master.address
			cpu_instruction_master_waitrequest                    => cpu_instruction_master_waitrequest,                        --                                                .waitrequest
			cpu_instruction_master_read                           => cpu_instruction_master_read,                               --                                                .read
			cpu_instruction_master_readdata                       => cpu_instruction_master_readdata,                           --                                                .readdata
			button_pio_s1_address                                 => mm_interconnect_0_button_pio_s1_address,                   --                                   button_pio_s1.address
			button_pio_s1_readdata                                => mm_interconnect_0_button_pio_s1_readdata,                  --                                                .readdata
			cpu_debug_mem_slave_address                           => mm_interconnect_0_cpu_debug_mem_slave_address,             --                             cpu_debug_mem_slave.address
			cpu_debug_mem_slave_write                             => mm_interconnect_0_cpu_debug_mem_slave_write,               --                                                .write
			cpu_debug_mem_slave_read                              => mm_interconnect_0_cpu_debug_mem_slave_read,                --                                                .read
			cpu_debug_mem_slave_readdata                          => mm_interconnect_0_cpu_debug_mem_slave_readdata,            --                                                .readdata
			cpu_debug_mem_slave_writedata                         => mm_interconnect_0_cpu_debug_mem_slave_writedata,           --                                                .writedata
			cpu_debug_mem_slave_byteenable                        => mm_interconnect_0_cpu_debug_mem_slave_byteenable,          --                                                .byteenable
			cpu_debug_mem_slave_waitrequest                       => mm_interconnect_0_cpu_debug_mem_slave_waitrequest,         --                                                .waitrequest
			cpu_debug_mem_slave_debugaccess                       => mm_interconnect_0_cpu_debug_mem_slave_debugaccess,         --                                                .debugaccess
			distance_in_s1_address                                => mm_interconnect_0_distance_in_s1_address,                  --                                  distance_in_s1.address
			distance_in_s1_readdata                               => mm_interconnect_0_distance_in_s1_readdata,                 --                                                .readdata
			jtag_uart_avalon_jtag_slave_address                   => mm_interconnect_0_jtag_uart_avalon_jtag_slave_address,     --                     jtag_uart_avalon_jtag_slave.address
			jtag_uart_avalon_jtag_slave_write                     => mm_interconnect_0_jtag_uart_avalon_jtag_slave_write,       --                                                .write
			jtag_uart_avalon_jtag_slave_read                      => mm_interconnect_0_jtag_uart_avalon_jtag_slave_read,        --                                                .read
			jtag_uart_avalon_jtag_slave_readdata                  => mm_interconnect_0_jtag_uart_avalon_jtag_slave_readdata,    --                                                .readdata
			jtag_uart_avalon_jtag_slave_writedata                 => mm_interconnect_0_jtag_uart_avalon_jtag_slave_writedata,   --                                                .writedata
			jtag_uart_avalon_jtag_slave_waitrequest               => mm_interconnect_0_jtag_uart_avalon_jtag_slave_waitrequest, --                                                .waitrequest
			jtag_uart_avalon_jtag_slave_chipselect                => mm_interconnect_0_jtag_uart_avalon_jtag_slave_chipselect,  --                                                .chipselect
			onchip_ram_s1_address                                 => mm_interconnect_0_onchip_ram_s1_address,                   --                                   onchip_ram_s1.address
			onchip_ram_s1_write                                   => mm_interconnect_0_onchip_ram_s1_write,                     --                                                .write
			onchip_ram_s1_readdata                                => mm_interconnect_0_onchip_ram_s1_readdata,                  --                                                .readdata
			onchip_ram_s1_writedata                               => mm_interconnect_0_onchip_ram_s1_writedata,                 --                                                .writedata
			onchip_ram_s1_byteenable                              => mm_interconnect_0_onchip_ram_s1_byteenable,                --                                                .byteenable
			onchip_ram_s1_chipselect                              => mm_interconnect_0_onchip_ram_s1_chipselect,                --                                                .chipselect
			onchip_ram_s1_clken                                   => mm_interconnect_0_onchip_ram_s1_clken,                     --                                                .clken
			pio_out_wd_s1_address                                 => mm_interconnect_0_pio_out_wd_s1_address,                   --                                   pio_out_wd_s1.address
			pio_out_wd_s1_write                                   => mm_interconnect_0_pio_out_wd_s1_write,                     --                                                .write
			pio_out_wd_s1_readdata                                => mm_interconnect_0_pio_out_wd_s1_readdata,                  --                                                .readdata
			pio_out_wd_s1_writedata                               => mm_interconnect_0_pio_out_wd_s1_writedata,                 --                                                .writedata
			pio_out_wd_s1_chipselect                              => mm_interconnect_0_pio_out_wd_s1_chipselect,                --                                                .chipselect
			pll_pll_slave_address                                 => mm_interconnect_0_pll_pll_slave_address,                   --                                   pll_pll_slave.address
			pll_pll_slave_write                                   => mm_interconnect_0_pll_pll_slave_write,                     --                                                .write
			pll_pll_slave_read                                    => mm_interconnect_0_pll_pll_slave_read,                      --                                                .read
			pll_pll_slave_readdata                                => mm_interconnect_0_pll_pll_slave_readdata,                  --                                                .readdata
			pll_pll_slave_writedata                               => mm_interconnect_0_pll_pll_slave_writedata,                 --                                                .writedata
			SERVO_HW_IP_0_avalon_slave_0_write                    => mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_write,      --                    SERVO_HW_IP_0_avalon_slave_0.write
			SERVO_HW_IP_0_avalon_slave_0_writedata                => mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_writedata,  --                                                .writedata
			SERVO_HW_IP_0_avalon_slave_0_chipselect               => mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_chipselect, --                                                .chipselect
			sierra_0_avalon_slave_0_address                       => mm_interconnect_0_sierra_0_avalon_slave_0_address,         --                         sierra_0_avalon_slave_0.address
			sierra_0_avalon_slave_0_write                         => mm_interconnect_0_sierra_0_avalon_slave_0_write,           --                                                .write
			sierra_0_avalon_slave_0_read                          => mm_interconnect_0_sierra_0_avalon_slave_0_read,            --                                                .read
			sierra_0_avalon_slave_0_readdata                      => mm_interconnect_0_sierra_0_avalon_slave_0_readdata,        --                                                .readdata
			sierra_0_avalon_slave_0_writedata                     => mm_interconnect_0_sierra_0_avalon_slave_0_writedata,       --                                                .writedata
			sierra_0_avalon_slave_0_chipselect                    => mm_interconnect_0_sierra_0_avalon_slave_0_chipselect,      --                                                .chipselect
			switch_pio_s1_address                                 => mm_interconnect_0_switch_pio_s1_address,                   --                                   switch_pio_s1.address
			switch_pio_s1_readdata                                => mm_interconnect_0_switch_pio_s1_readdata,                  --                                                .readdata
			sysid_control_slave_address                           => mm_interconnect_0_sysid_control_slave_address,             --                             sysid_control_slave.address
			sysid_control_slave_readdata                          => mm_interconnect_0_sysid_control_slave_readdata,            --                                                .readdata
			TIMER_HW_IP_0_avalon_slave_0_address                  => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_address,    --                    TIMER_HW_IP_0_avalon_slave_0.address
			TIMER_HW_IP_0_avalon_slave_0_write                    => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write,      --                                                .write
			TIMER_HW_IP_0_avalon_slave_0_read                     => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read,       --                                                .read
			TIMER_HW_IP_0_avalon_slave_0_readdata                 => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_readdata,   --                                                .readdata
			TIMER_HW_IP_0_avalon_slave_0_writedata                => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_writedata,  --                                                .writedata
			TIMER_HW_IP_0_avalon_slave_0_chipselect               => mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect, --                                                .chipselect
			VGA_IP_0_avalon_slave_0_address                       => mm_interconnect_0_vga_ip_0_avalon_slave_0_address,         --                         VGA_IP_0_avalon_slave_0.address
			VGA_IP_0_avalon_slave_0_write                         => mm_interconnect_0_vga_ip_0_avalon_slave_0_write,           --                                                .write
			VGA_IP_0_avalon_slave_0_read                          => mm_interconnect_0_vga_ip_0_avalon_slave_0_read,            --                                                .read
			VGA_IP_0_avalon_slave_0_readdata                      => mm_interconnect_0_vga_ip_0_avalon_slave_0_readdata,        --                                                .readdata
			VGA_IP_0_avalon_slave_0_writedata                     => mm_interconnect_0_vga_ip_0_avalon_slave_0_writedata,       --                                                .writedata
			VGA_IP_0_avalon_slave_0_chipselect                    => mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect       --                                                .chipselect
		);

	irq_mapper : component Range_finder_irq_mapper
		port map (
			clk           => pll_c0_clk,                     --       clk.clk
			reset         => rst_controller_reset_out_reset, -- clk_reset.reset
			receiver0_irq => irq_mapper_receiver0_irq,       -- receiver0.irq
			receiver1_irq => irq_mapper_receiver1_irq,       -- receiver1.irq
			sender_irq    => cpu_irq_irq                     --    sender.irq
		);

	rst_controller : component range_finder_rst_controller
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 1,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => pll_c0_clk,                         --       clk.clk
			reset_out      => rst_controller_reset_out_reset,     -- reset_out.reset
			reset_req      => rst_controller_reset_out_reset_req, --          .reset_req
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	rst_controller_001 : component range_finder_rst_controller_001
		generic map (
			NUM_RESET_INPUTS          => 2,
			OUTPUT_RESET_SYNC_EDGES   => "deassert",
			SYNC_DEPTH                => 2,
			RESET_REQUEST_PRESENT     => 0,
			RESET_REQ_WAIT_TIME       => 1,
			MIN_RST_ASSERTION_TIME    => 3,
			RESET_REQ_EARLY_DSRT_TIME => 1,
			USE_RESET_REQUEST_IN0     => 0,
			USE_RESET_REQUEST_IN1     => 0,
			USE_RESET_REQUEST_IN2     => 0,
			USE_RESET_REQUEST_IN3     => 0,
			USE_RESET_REQUEST_IN4     => 0,
			USE_RESET_REQUEST_IN5     => 0,
			USE_RESET_REQUEST_IN6     => 0,
			USE_RESET_REQUEST_IN7     => 0,
			USE_RESET_REQUEST_IN8     => 0,
			USE_RESET_REQUEST_IN9     => 0,
			USE_RESET_REQUEST_IN10    => 0,
			USE_RESET_REQUEST_IN11    => 0,
			USE_RESET_REQUEST_IN12    => 0,
			USE_RESET_REQUEST_IN13    => 0,
			USE_RESET_REQUEST_IN14    => 0,
			USE_RESET_REQUEST_IN15    => 0,
			ADAPT_RESET_REQUEST       => 0
		)
		port map (
			reset_in0      => reset_reset_n_ports_inv,            -- reset_in0.reset
			reset_in1      => cpu_debug_reset_request_reset,      -- reset_in1.reset
			clk            => clk_clk,                            --       clk.clk
			reset_out      => rst_controller_001_reset_out_reset, -- reset_out.reset
			reset_req      => open,                               -- (terminated)
			reset_req_in0  => '0',                                -- (terminated)
			reset_req_in1  => '0',                                -- (terminated)
			reset_in2      => '0',                                -- (terminated)
			reset_req_in2  => '0',                                -- (terminated)
			reset_in3      => '0',                                -- (terminated)
			reset_req_in3  => '0',                                -- (terminated)
			reset_in4      => '0',                                -- (terminated)
			reset_req_in4  => '0',                                -- (terminated)
			reset_in5      => '0',                                -- (terminated)
			reset_req_in5  => '0',                                -- (terminated)
			reset_in6      => '0',                                -- (terminated)
			reset_req_in6  => '0',                                -- (terminated)
			reset_in7      => '0',                                -- (terminated)
			reset_req_in7  => '0',                                -- (terminated)
			reset_in8      => '0',                                -- (terminated)
			reset_req_in8  => '0',                                -- (terminated)
			reset_in9      => '0',                                -- (terminated)
			reset_req_in9  => '0',                                -- (terminated)
			reset_in10     => '0',                                -- (terminated)
			reset_req_in10 => '0',                                -- (terminated)
			reset_in11     => '0',                                -- (terminated)
			reset_req_in11 => '0',                                -- (terminated)
			reset_in12     => '0',                                -- (terminated)
			reset_req_in12 => '0',                                -- (terminated)
			reset_in13     => '0',                                -- (terminated)
			reset_req_in13 => '0',                                -- (terminated)
			reset_in14     => '0',                                -- (terminated)
			reset_req_in14 => '0',                                -- (terminated)
			reset_in15     => '0',                                -- (terminated)
			reset_req_in15 => '0'                                 -- (terminated)
		);

	reset_reset_n_ports_inv <= not reset_reset_n;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_read_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_read;

	mm_interconnect_0_jtag_uart_avalon_jtag_slave_write_ports_inv <= not mm_interconnect_0_jtag_uart_avalon_jtag_slave_write;

	mm_interconnect_0_sierra_0_avalon_slave_0_chipselect_ports_inv <= not mm_interconnect_0_sierra_0_avalon_slave_0_chipselect;

	mm_interconnect_0_sierra_0_avalon_slave_0_read_ports_inv <= not mm_interconnect_0_sierra_0_avalon_slave_0_read;

	mm_interconnect_0_sierra_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_sierra_0_avalon_slave_0_write;

	mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect_ports_inv <= not mm_interconnect_0_vga_ip_0_avalon_slave_0_chipselect;

	mm_interconnect_0_vga_ip_0_avalon_slave_0_read_ports_inv <= not mm_interconnect_0_vga_ip_0_avalon_slave_0_read;

	mm_interconnect_0_vga_ip_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_vga_ip_0_avalon_slave_0_write;

	mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_chipselect_ports_inv <= not mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_chipselect;

	mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_servo_hw_ip_0_avalon_slave_0_write;

	mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect_ports_inv <= not mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_chipselect;

	mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read_ports_inv <= not mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_read;

	mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write_ports_inv <= not mm_interconnect_0_timer_hw_ip_0_avalon_slave_0_write;

	mm_interconnect_0_pio_out_wd_s1_write_ports_inv <= not mm_interconnect_0_pio_out_wd_s1_write;

	rst_controller_reset_out_reset_ports_inv <= not rst_controller_reset_out_reset;

end architecture rtl; -- of Range_finder
